module tt_um_riscv_core_top (
`ifdef USE_POWER_PINS
    input wire vccd1,   // 1.8V supply
    input wire vssd1,   // ground
`endif
    input  wire [7:0] ui_in,
    output wire [7:0] uo_out,
    input  wire [7:0] uio_in,
    output wire [7:0] uio_out,
    output wire [7:0] uio_oe,
    input  wire       ena,
    input  wire       clk,
    input  wire       rst_n
);


    // -------------------------------
    // GPIO REGISTER
    // -------------------------------
    wire [7:0] gpio_out;

    gpio_reg gpio_inst (
        .clk      (clk),
        .rst_n    (rst_n),
        .we       (uio_in[0] & ena),
        .wdata    (ui_in),
        .rdata    (),             // unused
        .gpio_out (gpio_out)
    );

    // -------------------------------
    // PWM GENERATOR
    // -------------------------------
    wire pwm_sig;

    pwm_generator pwm_inst (
        .clk     (clk),
        .rst_n   (rst_n),
        .duty    (gpio_out),
        .pwm_out (pwm_sig)
    );

    // -------------------------------
    // 7-SEG DISPLAY
    // -------------------------------
    wire [6:0] seg7;

    counter_to_7seg seg_inst (
        .val (gpio_out[3:0]),
        .seg (seg7)
    );

    // -------------------------------
    // OUTPUTS
    // -------------------------------
    assign uo_out  = gpio_out;
    assign uio_out = {pwm_sig, seg7};
    assign uio_oe  = 8'hFF;

endmodule
